package idma_proto_test;
  `include "idma_protocol_driver.sv"
  `include "idma_axi_driver.sv"
  `include "idma_source.sv"
endpackage : idma_proto_test